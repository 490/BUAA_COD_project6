`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:52:00 12/07/2014 
// Design Name: 
// Module Name:    gpr 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gpr(
    input Clk,
    input [4:0] A1,
    input [4:0] A2,
    input [4:0] A3,
    input We,
	 input Rst,
    input [31:0] WD,
    output [31:0] RD1,
    output [31:0] RD2
    );
/*=========================================================================================================*/
	reg [31:0] register[31:0];
/*=========================================================================================================*/
	integer i;
	initial
	begin
		for(i=0;i<33;i=i+1)
			register[i]<=32'b0;
	end
/*=========================================================================================================*/
	 always@(Rst)
	 begin
		for(i=0;i<=32;i=i+1)
			register[i]<=32'b0;
	 end
/*=========================================================================================================*/	
	//����ת��
	assign RD1=We?(A3==A1?(WD):(register[A1])):(register[A1]);
	assign RD2=We?(A3==A2?(WD):(register[A2])):(register[A2]);
/*=========================================================================================================*/
	always@(posedge Clk)
	begin
		if(We)
			register[A3]<=WD;
	end
/*=========================================================================================================*/
endmodule
