`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:53:47 12/07/2014 
// Design Name: 
// Module Name:    alu 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module alu(
    input [31:0] A,
    input [31:0] B,
    input [3:0] Op,
    output Over,
    output reg [31:0] C
    );
/*=========================================================================================================*/
	always@(*)
		begin
			case(Op[3:0])
				4'b0000:C=A+B;
				4'b0001:C=A-B;
				4'b0010:C=A|B;
				4'b0011:C=A&B;
				4'b0100:C=A^B;
				4'b0101:C=B<<(A%32);//sll,sllv
				4'b0110:C=B>>(A%32);//�߼�����srl
				4'b0111:			//��������sra							
							case(B[31])
								0:C=B>>(A%32);
								1:C=~(~B>>(A%32));
							endcase
				4'b1000:C=~(A|B);//nor
				4'b1001://�з���
							begin
							if(A>B) 
								C=32'b1;//С����1
							else
								C=0;//������0
							end
				4'b1010://�޷���
							begin
							if(A<B) 
								C=32'b1;//С����1
							else
								C=0;//������0
							end
							
			endcase
		end	
/*=========================================================================================================*/

/*=========================================================================================================*/
endmodule

